------------------------------
-- Elementos de Sistemas
-- Avaliacao Pratica 1
--
-- 10/2019
--
-- Questão 1
------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Questao1 is
  port (
	a : in  STD_LOGIC_VECTOR(2 downto 0);
	even : out STD_LOGIC := '0'	);
end entity;

architecture  rtl OF Questao1 IS

begin

end architecture;
