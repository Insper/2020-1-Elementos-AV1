------------------------------
-- Elementos de Sistemas
-- Avaliacao Pratica 1
--
-- 10/2019
--
-- Questão 5
------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Questao2 is
  port (
    x    : in  STD_LOGIC_VECTOR(1 downto 0);
    y    : in  STD_LOGIC_VECTOR(1 downto 0);
    xeqy : out STD_LOGIC;
    xlty : out STD_LOGIC);
end entity;

architecture  rtl OF Questao2 IS

begin


end architecture;
